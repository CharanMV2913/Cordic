/home/internals/Desktop/gpdk045_libfiles_1/gsclib045_tech.lef